// -----------------------------------------------------------------------------
// Universidade Federal do Recôncavo da Bahia
// -----------------------------------------------------------------------------
// Author : <seu nome aqui> <seu email>
// File   : DESim_top.sv
// Create : 2021-12-06 17:56:37
// Editor : Sublime Text 3, tab size (4)
// -----------------------------------------------------------------------------
// Module Purpose:
//    Top level interface from the DESim simulator
// -----------------------------------------------------------------------------
module top (
	////////////////////////	Clock Input	 	////////////////////////	 
	input wire CLOCK_50,
	////////////////////////	Push Button		////////////////////////
	input wire [3:0] KEY,
	////////////////////////	DPDT Switch		////////////////////////
	input wire 	[9:0] SW,
	////////////////////////	7-SEG Display   ////////////////////////
	output wire [6:0] HEX0
	);

	logic [3:0] digit;
	logic reset;

	//--------------------------------------------------------------------------
	assign digit = SW[3:0];
	assign reset = KEY[0];
	//--------------------------------------------------------------------------
	//	Output Logic
	//--------------------------------------------------------------------------
	dec7seg dec7seg_u0 ( 		,  		);
	//Instância do módulo hexto7seg
	//--------------------------------------------------------------------------	

endmodule
